
`timescale 1ns/1ps

module tb_MD5();

    reg i_Clk       ;
    reg i_Start     ;
    reg last512     ;
    reg i_Reset     ;
    reg [511:0] i_Data  ;

    wire[127:0] o_Data  ;
    wire o_FDone        ;
    wire o_FBusy        ;

MD5 md5(.i_clk(i_Clk),.i_start(i_Start),.last512(last512),.i_reset(i_Reset),.i_data(i_Data),.o_data(o_Data),.o_fBusy(o_FBusy),.o_fDone(o_FDone));

always #5i_Clk=~i_Clk;

initial begin
    i_Reset=1;
    i_Clk=1;
    i_Start=0;  
    last512=0;
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    i_Reset=0;  
    #20;
    i_Reset=1;
    #20;
    i_Start=1;  
    #10
    i_Start=0;  
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #10;
    i_Data=512'h61628000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_10000000_00000000; //ab
    #10;
    i_Data=512'h61626380_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_18000000_00000000; //abc
    #10;        
    i_Data=512'h61800000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_08000000_00000000; //a
    #800;
    last512=1;
    $stop;
end
endmodule